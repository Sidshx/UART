package uart_agent_pkg;
`include "uart_trans.sv"
`include "uart_gen.sv"
`include "uart_driver.sv"
`include "uart_monitor.sv"
`include "uart_agent.sv"

endpackage