package env_pkg;

import uart_agent_pkg::*;
`include "uart_scoreboard.sv"
`include "env.sv"

endpackage
